magic
tech scmos
timestamp 1550265184
<< nwell >>
rect 0 -4 24 25
rect 30 -4 86 25
rect 92 -4 164 25
rect 170 -4 194 25
<< ntransistor >>
rect 11 -24 13 -20
rect 181 -17 183 -13
rect 41 -43 43 -39
rect 49 -43 51 -39
rect 57 -43 59 -39
rect 65 -43 67 -39
rect 73 -43 75 -39
rect 103 -43 105 -39
rect 111 -43 113 -39
rect 119 -43 121 -39
rect 127 -43 129 -39
rect 135 -43 137 -39
rect 143 -43 145 -39
rect 151 -43 153 -39
<< ptransistor >>
rect 11 2 13 14
rect 41 2 43 14
rect 49 2 51 14
rect 57 2 59 14
rect 65 2 67 14
rect 73 2 75 14
rect 103 2 105 14
rect 111 2 113 14
rect 119 2 121 14
rect 127 2 129 14
rect 135 2 137 14
rect 143 2 145 14
rect 151 2 153 14
rect 181 2 183 14
<< ndiffusion >>
rect 10 -24 11 -20
rect 13 -24 14 -20
rect 180 -17 181 -13
rect 183 -17 184 -13
rect 40 -43 41 -39
rect 43 -43 44 -39
rect 48 -43 49 -39
rect 51 -43 52 -39
rect 56 -43 57 -39
rect 59 -43 60 -39
rect 64 -43 65 -39
rect 67 -43 73 -39
rect 75 -43 76 -39
rect 102 -43 103 -39
rect 105 -43 111 -39
rect 113 -43 119 -39
rect 121 -43 122 -39
rect 126 -43 127 -39
rect 129 -43 130 -39
rect 134 -43 135 -39
rect 137 -43 138 -39
rect 142 -43 143 -39
rect 145 -43 146 -39
rect 150 -43 151 -39
rect 153 -43 154 -39
<< pdiffusion >>
rect 10 2 11 14
rect 13 2 14 14
rect 40 2 41 14
rect 43 2 49 14
rect 51 2 52 14
rect 56 2 57 14
rect 59 2 60 14
rect 64 2 65 14
rect 67 2 68 14
rect 72 2 73 14
rect 75 2 76 14
rect 102 2 103 14
rect 105 2 106 14
rect 110 2 111 14
rect 113 2 114 14
rect 118 2 119 14
rect 121 2 122 14
rect 126 2 127 14
rect 129 2 135 14
rect 137 2 143 14
rect 145 2 146 14
rect 150 2 151 14
rect 153 2 154 14
rect 180 2 181 14
rect 183 2 184 14
<< ndcontact >>
rect 6 -24 10 -20
rect 14 -24 18 -20
rect 176 -17 180 -13
rect 184 -17 188 -13
rect 36 -43 40 -39
rect 44 -43 48 -39
rect 52 -43 56 -39
rect 60 -43 64 -39
rect 76 -43 80 -39
rect 98 -43 102 -39
rect 122 -43 126 -39
rect 130 -43 134 -39
rect 138 -43 142 -39
rect 146 -43 150 -39
rect 154 -43 158 -39
<< pdcontact >>
rect 6 2 10 14
rect 14 2 18 14
rect 36 2 40 14
rect 52 2 56 14
rect 60 2 64 14
rect 68 2 72 14
rect 76 2 80 14
rect 98 2 102 14
rect 106 2 110 14
rect 114 2 118 14
rect 122 2 126 14
rect 146 2 150 14
rect 154 2 158 14
rect 176 2 180 14
rect 184 2 188 14
<< psubstratepcontact >>
rect 14 -46 18 -42
rect 88 -46 92 -42
rect 176 -46 180 -42
<< nsubstratencontact >>
rect 14 18 18 22
rect 68 18 72 22
rect 98 18 102 22
rect 114 18 118 22
rect 176 18 180 22
<< polysilicon >>
rect 11 14 13 16
rect 41 14 43 16
rect 49 14 51 16
rect 57 14 59 16
rect 65 14 67 16
rect 73 14 75 16
rect 103 14 105 16
rect 111 14 113 16
rect 119 14 121 16
rect 127 14 129 16
rect 135 14 137 16
rect 143 14 145 16
rect 151 14 153 16
rect 181 14 183 16
rect 11 -20 13 2
rect 41 -20 43 2
rect 11 -26 13 -24
rect 41 -39 43 -24
rect 49 -26 51 2
rect 57 -13 59 2
rect 49 -39 51 -30
rect 57 -39 59 -17
rect 65 -19 67 2
rect 65 -39 67 -23
rect 73 -26 75 2
rect 103 -19 105 2
rect 73 -39 75 -30
rect 103 -39 105 -23
rect 111 -26 113 2
rect 119 -13 121 2
rect 111 -39 113 -30
rect 119 -39 121 -17
rect 127 -19 129 2
rect 127 -39 129 -23
rect 135 -25 137 2
rect 143 -13 145 2
rect 151 -7 153 2
rect 135 -39 137 -29
rect 143 -39 145 -17
rect 151 -39 153 -11
rect 181 -13 183 2
rect 181 -19 183 -17
rect 41 -45 43 -43
rect 49 -45 51 -43
rect 57 -45 59 -43
rect 65 -45 67 -43
rect 73 -45 75 -43
rect 103 -45 105 -43
rect 111 -45 113 -43
rect 119 -45 121 -43
rect 127 -45 129 -43
rect 135 -45 137 -43
rect 143 -45 145 -43
rect 151 -45 153 -43
<< polycontact >>
rect 13 -10 17 -6
rect 40 -24 44 -20
rect 56 -17 60 -13
rect 48 -30 52 -26
rect 64 -23 68 -19
rect 102 -23 106 -19
rect 72 -30 76 -26
rect 118 -17 122 -13
rect 110 -30 114 -26
rect 126 -23 130 -19
rect 177 -5 181 -1
rect 150 -11 154 -7
rect 142 -17 146 -13
rect 134 -29 138 -25
<< metal1 >>
rect 0 23 194 27
rect 14 22 18 23
rect 68 22 72 23
rect 14 14 18 18
rect 36 17 64 20
rect 36 14 40 17
rect 60 14 64 17
rect 6 -20 10 2
rect 52 -7 56 2
rect 68 14 72 18
rect 98 22 102 23
rect 98 14 102 18
rect 114 22 118 23
rect 176 22 180 23
rect 114 14 118 18
rect 122 17 158 20
rect 122 14 126 17
rect 154 14 158 17
rect 60 -1 64 2
rect 76 -1 80 2
rect 60 -4 80 -1
rect 106 -1 110 2
rect 122 -1 126 2
rect 106 -4 126 -1
rect 176 14 180 18
rect 146 -1 150 2
rect 146 -4 177 -1
rect 17 -10 150 -7
rect 14 -42 18 -24
rect 28 -32 32 -10
rect 60 -16 87 -13
rect 91 -16 118 -13
rect 122 -16 142 -13
rect 44 -23 64 -20
rect 68 -23 102 -20
rect 106 -23 126 -20
rect 52 -29 72 -26
rect 76 -29 110 -26
rect 114 -29 134 -26
rect 161 -32 165 -4
rect 184 -13 188 2
rect 36 -36 56 -33
rect 36 -39 40 -36
rect 52 -39 56 -36
rect 60 -39 64 -36
rect 98 -39 102 -36
rect 130 -36 150 -33
rect 130 -39 134 -36
rect 146 -39 150 -36
rect 44 -46 48 -43
rect 76 -46 80 -43
rect 158 -36 165 -32
rect 154 -39 158 -36
rect 176 -42 180 -17
rect 122 -46 126 -43
rect 138 -46 142 -43
rect 0 -50 194 -46
<< m2contact >>
rect 87 -17 91 -13
rect 28 -36 32 -32
rect 60 -36 64 -32
rect 98 -36 102 -32
rect 154 -36 158 -32
<< metal2 >>
rect 32 -36 60 -32
rect 102 -36 154 -32
<< labels >>
rlabel metal1 8 -7 8 -7 1 COUT
rlabel metal1 89 25 89 25 5 vdd
rlabel metal1 90 -48 90 -48 1 gnd
rlabel metal1 186 -7 186 -7 1 SUM
rlabel polycontact 50 -28 50 -28 1 B
rlabel polycontact 58 -15 58 -15 1 CIN
rlabel polycontact 42 -22 42 -22 1 A
<< end >>
